module not_4(out,in);
	input[3:0] in;
	output[3:0] out;
	not not1(out[0],in[0]);
	not not2(out[1],in[1]);
	not not3(out[2],in[2]);
	not not4(out[3],in[3]);
endmodule
	