/*module FSM_buf(in,Current_state,New_state);
	input[2:0] Current_state;
	input in;
	output out;
	//if (in==1'b1)
	 //New_state=(Current_state+1)/4;
endmodule
*/